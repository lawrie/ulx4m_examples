module top (
    output [3:0] led
);
    assign led = 4'b1001;

endmodule
